module resource

import mv.thirdparty.cute as sb

pub struct Spritebatcher {
pub mut:
	config   sb.SpritebatchConfig
	batcher  ?sb.Spritebatch
	textures []&Texture
}
