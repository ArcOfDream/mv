module math

pub enum Axis {
	x
	y
}
