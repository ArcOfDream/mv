module resource

pub struct RresFile {
pub:
	resource_type ResourceType = .archive
pub mut:
	name string
}
