module util
