module util

// import vres
// import mv.resource as r

// pub fn unpack_resource_chunk(chunk &vres.ResourceChunk) {}

// pub fn load_texture_from_resource_chunk(chunk &vres.ResourceChunk) ?r.Texture {
// 	if chunk.info.compType == .rres_comp_none && chunk.info.cipherType == .rres_cipher_none {

// 	}

// 	return r.Texture{}
// }
